


"Title:unknown_tag"
Footage of a Ukrainian FPV drone intercepting a Russian UAV flying a Soviet victory banner.
Timestamp: 3:40 AM · Jun 3, 2025
--Footage_of_a_Ukrainian_FPV_drone_intercepting_a_Russian_UAV_image_1_143831.jpg
--Footage_of_a_Ukrainian_FPV_drone_intercepting_a_Russian_UAV_143832.mp4
https://x.com/Osinttechnical/status/1929624125632643187

cc-Source- https://t.me/robert_magyar/1115… | Additional footage of Magyar’s unit downing dozens of Russian fixed wing drones.
cc-That banner would make one helluva souvenir  | (or ass-wipe )
cc-DE PAUVRE POMER SOVIÉTIQUE ... apart joué aux GUIGNOLS c'est tout ce qu ils peuvent avoir comme exploits... Les jours ont compté de maintenant signer leurs FIN MONDIALE.
cc-Based
cc-Fully missed it
cc-NSW’s State of Origin squad has been rocked by injury carnage, while the Maroons are set to blood a shock bolter in the series opener.


"Title:unknown_tag"
Norway will help Ukraine cover a potential one billion euro ($1.08 billion) gas deficit, President Volodymyr Zelensky announced following a meeting with Norwegian Prime Minister Jonas Gahr Store in Vilnius on June 2.
Timestamp: 7:37 AM · Jun 3, 2025
https://x.com/KyivIndependent/status/1929683748372860933

cc-Better Norway than us.  Thanks Norway!
cc-This isn’t the American families problem
cc-The truth behind the shotgun.  This story changed my life. I hope it can help you. Read the first couple of chapters for free on Amazon: https://mybook.to/oBjJGA?twclid=27b4hlkx8mia1dwfxtwvdincu7
cc-Ukraine is nothing more than a rump state at this point. Taking handouts from the entire world. Sad
cc-Nice
cc-Solidarity means nurturing reciprocal relationships. Trumps America is about exploiting those kinds of relationships The Norwegians like most of Europe's Union partners know why Solidarity is so important.  | What a great example to Americans. Currently, we're stuck in a me world


"Title:unknown_tag"
Typhoon Cremee Trucks
Timestamp: 5:37 AM · Jun 3, 2025
--Typhoon_Cremee_Trucks_image_1_143852.jpg
--Typhoon_Cremee_Trucks_image_2_143853.jpg
https://x.com/Schizointel/status/1929668709263855883


   "Quoted Tweet:"

Again, no one would mistake a 150 ft long, olive-drab Typhon launcher that has a gross combined weight rating in excess of 70 tons with ... a civilian Mister Softee truck.
Timestamp: 5:35 AM · Jun 3, 2025
--Again_no_one_would_mistake_a_150_ft_long_olive-drab_image_1_143901.jpg
--Again_no_one_would_mistake_a_150_ft_long_olive-drab_image_2_143902.jpg
https://x.com/ArmsControlWonk/status/1929653621685416380


   "Quoted Tweet:"

cc-Russia literally exports cruise missiles disguised as shipping containers.
cc-The US too. | Behold, from 2023...
cc-Exactly


"Title:unknown_tag"
Images of reportedly the power station near  occupied Melitopol that was hit and is now ablaze. Power has been knocked out in the area.
Timestamp: 4:57 AM · Jun 3, 2025
--Images_of_reportedly_the_power_station_near_occupied_Melitopol_th_image_1_143918.jpg
--Images_of_reportedly_the_power_station_near_occupied_Melitopol_th_image_2_143919.jpg
--Images_of_reportedly_the_power_station_near_occupied_Melitopol_th_image_3_143920.jpg
--Images_of_reportedly_the_power_station_near_occupied_Melitopol_th_image_4_143921.jpg
https://x.com/raging545/status/1929643602139058193

cc-pic 2/4 | Purported fire at  Electrical Substation Melitopol   | PoV ~ 46.839138, 35.352841 | @GeoConfirmed |  @UAControlMap |  @giK1893


"Title:unknown_tag"
It’s Not a Tiny House—It’s Ukrainian FPV Drone Launcher

The containers look like tiny homes—solar panels on top, an empty interior, nothing suspicious. 

But inside, they charge batteries and hide a drone just 20 cm below the ceiling.

Even if you step in, you wouldn’t notice it. The roof opens using a motorized rail or belt.
A weak corner bracket breaks under pressure, dropping the roof.
As the motor keeps running, it forces the roof open and ejects it.
The falling roof hits the side wall—proof it opens and drops in one motion.

A stealthy drone launch system, disguised as a harmless cabin.
Timestamp: 3:35 AM · Jun 3, 2025
--Its_Not_a_Tiny_HouseIts_Ukrainian_FPV_Drone_Launcher_The_image_1_143931.jpg
--Its_Not_a_Tiny_HouseIts_Ukrainian_FPV_Drone_Launcher_The_image_2_143931.jpg
--Its_Not_a_Tiny_HouseIts_Ukrainian_FPV_Drone_Launcher_The_image_3_143932.jpg
--Its_Not_a_Tiny_HouseIts_Ukrainian_FPV_Drone_Launcher_The_image_4_143932.jpg
https://x.com/clashreport/status/1929622853462512000

cc-これはタイニーハウスではありません。ウクライナのFPVドローンランチャーです。 | コンテナは小さな家のように見えます。上にはソーラーパネルがあり、内部は空っぽで、何も不審な点はありません。 | しかし、内部ではバッテリーを充電し、天井からわずか20センチ下にドローンを隠しています。
cc-I dont support Ukraine, but this was genius
cc-After some time, Ukranians will hunt for the man who came up with the idea. #RussiaUkraineWar #Russia
cc-The truth behind the shotgun.  This story changed my life. I hope it can help you. Read the first couple of chapters for free on Amazon: https://mybook.to/oBjJGA?twclid=2vrk80ppwckmpdjjky53pv2hm
cc-Geee...wonder where they got the idea
cc-@CedricLeighton |  perfect disguise - a shipping container painted any scheme or distressed to hide it's age.....portable morgue?


"Title:unknown_tag"
Zelensky says he's ready to meet with Putin, Trump in Turkey. 

"I told (Turkish President) that I support a meeting at the level of leaders, because I have the impression that there will be no ceasefire without our meeting," Zelensky said on June 2.
Timestamp: 6:06 AM · Jun 3, 2025
https://x.com/KyivIndependent/status/1929660852250329412

cc-Representation from European leaders is essential.
cc-
cc-Canadian-born new Greens leader Larissa Waters made headlines in 2017 for one infamous Parliament act.
cc-putler won't go to Turkey, as there exists no bunkers equivalent to the one at home
cc-I'm becoming rather eclectic about a peaceful solution.
cc-pootie will avoid that meeting like the plague.


"Title:unknown_tag"
Massive drones attack on Crimea 

Map from 
@DrnBmbr
Timestamp: 4:49 AM · Jun 3, 2025
--Massive_drones_attack_on_Crimea_Map_from_DrnBmbr_image_1_144005.jpg
https://x.com/Maks_NAFO_FELLA/status/1929641637002592568

cc-Overload the bridge air defense with drones and then send in the ballistics, Taurus, and Storm Shadows.
cc-Weren't the remains of the Black Sea Fleet moved to Eastern Crimea?
cc-The truth behind the shotgun.  This story changed my life. I hope it can help you. Read the first couple of chapters for free on Amazon: https://mybook.to/oBjJGA?twclid=24f36ghsh6g43nmq4um0pt02qc
cc-On eastern Crimea ...
cc-Holy fuck
cc-How does Dronbomber get this info? These are really good products but how legit are they?


"Title:unknown_tag"
Melitopol is completely without power.
Timestamp: 4:19 AM · Jun 3, 2025
--Melitopol_is_completely_without_power_image_1_144014.jpg
https://x.com/Maks_NAFO_FELLA/status/1929634067882148227

cc-Things are happening...
cc-UKRAINE strikes of RUSSIAN strikes!!
cc-Access global liquidity. Tighter spreads. T+0 settlements. Personalised service.
cc-Melitopol is completely without power (including cell towers) | If one wanted to hide approach of drones or Taurus missiles on oproach to Kerch Bridge, it would make sense to cut power to occupied areas that might otherwise warn others...


"Title:unknown_tag"
Occupied Melitopol… BAVOVNA 
Timestamp: 4:00 AM · Jun 3, 2025
--Occupied_Melitopol_BAVOVNA_image_1_144024.jpg
https://x.com/Maks_NAFO_FELLA/status/1929629266473255249

cc-Ocrs
cc-I BAVOVNA looks flaming lovely
cc-Feminists are HURTING Women and Men By Pushing their Sexist Man-hatred in the domestic violence crisis.  Hijacking a tragic and important issue for their own sick political gain.   | It’s time brave men all stood up and called it out.   I’ll start…
cc-Melitopol is Ukraine
cc-Bavovna!


"Title:unknown_tag"
The Russian delegation is not as cheerful as in the past negotiations with Ukraine.
Timestamp: 8:02 PM · Jun 2, 2025
--The_Russian_delegation_is_not_as_cheerful_as_in_the_image_1_144045.jpg
--The_Russian_delegation_is_not_as_cheerful_as_in_the_144046.mp4
https://x.com/Maks_NAFO_FELLA/status/1929509020907253936

cc-None of them have a choice or power to make a Decision lol
cc-They are not interested in negotiations!
cc-Trade crypto on the go with the BTC Markets mobile app.
cc-How did they arrive at these "negotiations" ? If it was by aircraft, is it where they left it?
cc-Ukraine should have brought some toy trucks to put on their table.
cc-Their scare of falling out of windows. | I bet they asked for all the windows to be close before they started negotiating.


"Title:unknown_tag"
85 hours left
Timestamp: 5:31 AM · Jun 3, 2025
--85_hours_left_image_1_144058.jpg
--85_hours_left_144059.mp4
https://x.com/Prune602/status/1929652222704357487

cc-83.....
cc-80 hrs 54 minutes
cc-I would be suprised by another key rate increase at this point. To me it looks as if Kremlin has given out the order to Central Bank to not worsen the credit situation. They cannot stop inflation this way anyways as long as Kremlin throws out money left and right. But lets see
cc-Discover the software trusted by home building professionals: architects, builders, designers, and lumberyards all agree that SoftPlan is the top choice for drawing houses.
cc-Didn’t Putin say that they are not  allowed to raise it.


"Title:unknown_tag"
Ukraine's largest private energy company DTEK secured a $72-million loan to build one of the largest battery energy storage complexes in Eastern Europe, the company said on June 3.
Timestamp: 5:22 AM · Jun 3, 2025
https://x.com/KyivIndependent/status/1929649753757044784

cc-* | Yet another inorganic U.S  | Taxpayer funded foreign aid business venture.  | Social Welfare...for Ukraine
cc-Anybody who lends money for this needs to have his head examined (or be investigate for fraud). | Nearly 100% probability it will get destroyed.
cc-Awesome!!!!!
cc-Great project, but why now? You just know Russia will just destroy it and it will become a waste of $72 million.
cc-Decentralize them Ukraine, so they can’t be blown up! Put a battery in every building.
cc-ukraine investing in energy storage is smart. it’s about reducing dependence on moscovite energy, boosting our resilience, and building a real economy. no more reliance on moscovite cash flows. we keep fighting, we keep building.


"Title:unknown_tag"
Russia is in real trouble. Western sanctions have cut daily seaborne oil exports from 4 million barrels per day in January 2025 to 3 million now. This is before UK and EU sanctions - announced this month - have even fully hit. Putin's money machine is under real pressure now...
Timestamp: 3:32 PM · May 30, 2025
--Russia_is_in_real_trouble_Western_sanctions_have_cut_daily_image_1_144121.jpg
https://x.com/robin_j_brooks/status/1928353917714211031

cc-Wow look at this - Greece should be ashamed of themselves...
cc-Any nations still buying KGB Putin's energy (natural gas/crude oil) via his fleet of ghost supertankers should be hit with stiff import duty fees on their exports.
cc-Can you provide a chart of yourself, number of hours day dreaming?
cc-WIN the ultimate State of Origin Game 3 experience!  | Prize includes: |  2 x diamond passes to Origin Game 3 on the 9th July, 2025 |  2 nights at the Pullman Olympic park with breakfast & late check out (9-11th July) |  $1,500AUD Prezzee Smart eGift card to use towards flights
cc-To bad we have a russia shill in the WH
cc-Should have been done when they invaded ukraine.


"Title:unknown_tag"
Melitpol is reportedly completely out of power after Ukrainian drone attacks.
Timestamp: 4:06 AM · Jun 3, 2025
--Melitpol_is_reportedly_completely_out_of_power_after_Ukrainian_dr_image_1_144149.jpg
--Melitpol_is_reportedly_completely_out_of_power_after_Ukrainian_dr_image_2_144150.jpg
https://x.com/NOELreports/status/1929638659726127596


   "Quoted Tweet:"

Timestamp: 4:06 AM · Jun 3, 2025
--Reports_indicate_a_large_wave_of_Ukrainian_drones_flying_over_image_1_144157.jpg
https://x.com/NOELreports/status/1929630752217645074

cc-Reports indicate a large wave of Ukrainian drones flying over occupied Enerhodar and Berdiansk, heading toward occupied Crimea and the Kuban region.
cc-In occupied Melitopol, explosions were reported and parts of the city are without power.
cc-ukraine’s drone game isn’t just about hitting targets — it’s about showing moscovia they’re losing ground everywhere, even in their own backyard. night missions like this keep their illusions of control shattered. they can’t hide from our tech.
cc-You are not just a dog, you are my sanity, my happiness, my teacher, my therapist and my best friend   | Get it https://warmwishmall.co/dog-craft?twclid=2-5jyeay9qy7cnd2vjrgcz30png
cc-




"Title:unknown_tag"

--Melitpol_is_reportedly_completely_out_of_power_after_Ukrainian_dr_image_1_144149.jpg
--Melitpol_is_reportedly_completely_out_of_power_after_Ukrainian_dr_image_2_144150.jpg
https://x.com/NOELreports/status/1929638659726127596


   "Quoted Tweet:"

Reports indicate a large wave of Ukrainian drones flying over occupied Enerhodar and Berdiansk, heading toward occupied Crimea and the Kuban region.
Timestamp: 4:06 AM · Jun 3, 2025
--Reports_indicate_a_large_wave_of_Ukrainian_drones_flying_over_image_1_144157.jpg
https://x.com/NOELreports/status/1929630752217645074

cc-Reports indicate a large wave of Ukrainian drones flying over occupied Enerhodar and Berdiansk, heading toward occupied Crimea and the Kuban region.
cc-In occupied Melitopol, explosions were reported and parts of the city are without power.
cc-ukraine’s drone game isn’t just about hitting targets — it’s about showing moscovia they’re losing ground everywhere, even in their own backyard. night missions like this keep their illusions of control shattered. they can’t hide from our tech.
cc-You are not just a dog, you are my sanity, my happiness, my teacher, my therapist and my best friend   | Get it https://warmwishmall.co/dog-craft?twclid=2-5jyeay9qy7cnd2vjrgcz30png
cc-

