


"Title:unknown_tag"
Footage of a Ukrainian FPV drone intercepting a Russian UAV flying a Soviet victory banner.




"Title:unknown_tag"
Norway will help Ukraine cover a potential one billion euro ($1.08 billion) gas deficit, President Volodymyr Zelensky announced following a meeting with Norwegian Prime Minister Jonas Gahr Store in Vilnius on June 2.




"Title:unknown_tag"
Typhoon Cremee Trucks




"Title:unknown_tag"
Images of reportedly the power station near  occupied Melitopol that was hit and is now ablaze. Power has been knocked out in the area.




"Title:unknown_tag"
It’s Not a Tiny House—It’s Ukrainian FPV Drone Launcher




"Title:unknown_tag"
Zelensky says he's ready to meet with Putin, Trump in Turkey. 




"Title:unknown_tag"
Massive drones attack on Crimea 
Melitopol is completely without power.




"Title:unknown_tag"
Occupied Melitopol… BAVOVNA 




"Title:unknown_tag"
The Russian delegation is not as cheerful as in the past negotiations with Ukraine.




"Title:unknown_tag"
85 hours left




"Title:unknown_tag"
Ukraine's largest private energy company DTEK secured a $72-million loan to build one of the largest battery energy storage complexes in Eastern Europe, the company said on June 3.

"Title:Economy"

Russia is in real trouble. Western sanctions have cut daily seaborne oil exports from 4 million barrels per day in January 2025 to 3 million now. This is before UK and EU sanctions - announced this month - have even fully hit. Putin's money machine is under real pressure now...

"Title:Politics"

"Title:Part3"

"Title:Part4"




"Title:unknown_tag"
Melitpol is reportedly completely out of power after Ukrainian drone attacks.